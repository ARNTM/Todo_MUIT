module top();
      nios_system_tb tb ();
      test_program pgm ();
endmodule
