
module nios_system (
	clk_50_in_clk,
	reset_reset_n);	

	input		clk_50_in_clk;
	input		reset_reset_n;
endmodule
