// nios_system.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module nios_system (
		input  wire  clk_50_in_clk, // clk_50_in.clk
		input  wire  reset_reset_n  //     reset.reset_n
	);

	wire  [31:0] mm_master_bfm_m0_readdata;                                 // mm_interconnect_0:mm_master_bfm_m0_readdata -> mm_master_bfm:avm_readdata
	wire         mm_master_bfm_m0_waitrequest;                              // mm_interconnect_0:mm_master_bfm_m0_waitrequest -> mm_master_bfm:avm_waitrequest
	wire   [2:0] mm_master_bfm_m0_address;                                  // mm_master_bfm:avm_address -> mm_interconnect_0:mm_master_bfm_m0_address
	wire         mm_master_bfm_m0_read;                                     // mm_master_bfm:avm_read -> mm_interconnect_0:mm_master_bfm_m0_read
	wire  [31:0] mm_master_bfm_m0_writedata;                                // mm_master_bfm:avm_writedata -> mm_interconnect_0:mm_master_bfm_m0_writedata
	wire         mm_master_bfm_m0_write;                                    // mm_master_bfm:avm_write -> mm_interconnect_0:mm_master_bfm_m0_write
	wire         mm_interconnect_0_chromaprocessor_avalon_slave_chipselect; // mm_interconnect_0:ChromaProcessor_avalon_slave_chipselect -> ChromaProcessor:chipselect
	wire  [31:0] mm_interconnect_0_chromaprocessor_avalon_slave_readdata;   // ChromaProcessor:readdata -> mm_interconnect_0:ChromaProcessor_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_chromaprocessor_avalon_slave_address;    // mm_interconnect_0:ChromaProcessor_avalon_slave_address -> ChromaProcessor:address
	wire         mm_interconnect_0_chromaprocessor_avalon_slave_read;       // mm_interconnect_0:ChromaProcessor_avalon_slave_read -> ChromaProcessor:read
	wire         mm_interconnect_0_chromaprocessor_avalon_slave_write;      // mm_interconnect_0:ChromaProcessor_avalon_slave_write -> ChromaProcessor:write
	wire  [31:0] mm_interconnect_0_chromaprocessor_avalon_slave_writedata;  // mm_interconnect_0:ChromaProcessor_avalon_slave_writedata -> ChromaProcessor:writedata
	wire         chromaprocessor_avalon_streaming_source_valid;             // ChromaProcessor:output_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] chromaprocessor_avalon_streaming_source_data;              // ChromaProcessor:output_data -> avalon_st_adapter:in_0_data
	wire         chromaprocessor_avalon_streaming_source_ready;             // avalon_st_adapter:in_0_ready -> ChromaProcessor:output_ready
	wire         chromaprocessor_avalon_streaming_source_startofpacket;     // ChromaProcessor:output_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         chromaprocessor_avalon_streaming_source_endofpacket;       // ChromaProcessor:output_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire   [1:0] chromaprocessor_avalon_streaming_source_empty;             // ChromaProcessor:output_empty -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                             // avalon_st_adapter:out_0_valid -> st_sink_bfm:sink_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                              // avalon_st_adapter:out_0_data -> st_sink_bfm:sink_data
	wire         avalon_st_adapter_out_0_ready;                             // st_sink_bfm:sink_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                     // avalon_st_adapter:out_0_startofpacket -> st_sink_bfm:sink_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                       // avalon_st_adapter:out_0_endofpacket -> st_sink_bfm:sink_endofpacket
	wire   [0:0] st_source_bfm_background_src_valid;                        // st_source_bfm_background:src_valid -> avalon_st_adapter_001:in_0_valid
	wire  [29:0] st_source_bfm_background_src_data;                         // st_source_bfm_background:src_data -> avalon_st_adapter_001:in_0_data
	wire         st_source_bfm_background_src_ready;                        // avalon_st_adapter_001:in_0_ready -> st_source_bfm_background:src_ready
	wire   [0:0] st_source_bfm_background_src_startofpacket;                // st_source_bfm_background:src_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire   [0:0] st_source_bfm_background_src_endofpacket;                  // st_source_bfm_background:src_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;                         // avalon_st_adapter_001:out_0_valid -> ChromaProcessor:pixel_fondo_valid
	wire  [29:0] avalon_st_adapter_001_out_0_data;                          // avalon_st_adapter_001:out_0_data -> ChromaProcessor:pixel_fondo
	wire         avalon_st_adapter_001_out_0_ready;                         // ChromaProcessor:pixel_fondo_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;                 // avalon_st_adapter_001:out_0_startofpacket -> ChromaProcessor:pixel_fondo_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                   // avalon_st_adapter_001:out_0_endofpacket -> ChromaProcessor:pixel_fondo_endofpacket
	wire   [1:0] avalon_st_adapter_001_out_0_empty;                         // avalon_st_adapter_001:out_0_empty -> ChromaProcessor:pixel_fondo_empty
	wire   [0:0] st_source_bfm_foreground_src_valid;                        // st_source_bfm_foreground:src_valid -> avalon_st_adapter_002:in_0_valid
	wire  [29:0] st_source_bfm_foreground_src_data;                         // st_source_bfm_foreground:src_data -> avalon_st_adapter_002:in_0_data
	wire         st_source_bfm_foreground_src_ready;                        // avalon_st_adapter_002:in_0_ready -> st_source_bfm_foreground:src_ready
	wire   [0:0] st_source_bfm_foreground_src_startofpacket;                // st_source_bfm_foreground:src_startofpacket -> avalon_st_adapter_002:in_0_startofpacket
	wire   [0:0] st_source_bfm_foreground_src_endofpacket;                  // st_source_bfm_foreground:src_endofpacket -> avalon_st_adapter_002:in_0_endofpacket
	wire         avalon_st_adapter_002_out_0_valid;                         // avalon_st_adapter_002:out_0_valid -> ChromaProcessor:pixel_video_valid
	wire  [29:0] avalon_st_adapter_002_out_0_data;                          // avalon_st_adapter_002:out_0_data -> ChromaProcessor:pixel_video
	wire         avalon_st_adapter_002_out_0_ready;                         // ChromaProcessor:pixel_video_ready -> avalon_st_adapter_002:out_0_ready
	wire         avalon_st_adapter_002_out_0_startofpacket;                 // avalon_st_adapter_002:out_0_startofpacket -> ChromaProcessor:pixel_video_startofpacket
	wire         avalon_st_adapter_002_out_0_endofpacket;                   // avalon_st_adapter_002:out_0_endofpacket -> ChromaProcessor:pixel_video_endofpacket
	wire   [1:0] avalon_st_adapter_002_out_0_empty;                         // avalon_st_adapter_002:out_0_empty -> ChromaProcessor:pixel_video_empty
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [ChromaProcessor:reset, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, mm_interconnect_0:mm_master_bfm_clk_reset_reset_bridge_in_reset_reset, mm_master_bfm:reset, st_sink_bfm:reset, st_source_bfm_background:reset, st_source_bfm_foreground:reset]

	altera_up_avalon_chroma_key chromaprocessor (
		.clk                       (clk_50_in_clk),                                             //                   clock.clk
		.reset                     (rst_controller_reset_out_reset),                            //                   reset.reset
		.output_data               (chromaprocessor_avalon_streaming_source_data),              // avalon_streaming_source.data
		.output_empty              (chromaprocessor_avalon_streaming_source_empty),             //                        .empty
		.output_ready              (chromaprocessor_avalon_streaming_source_ready),             //                        .ready
		.output_startofpacket      (chromaprocessor_avalon_streaming_source_startofpacket),     //                        .startofpacket
		.output_valid              (chromaprocessor_avalon_streaming_source_valid),             //                        .valid
		.output_endofpacket        (chromaprocessor_avalon_streaming_source_endofpacket),       //                        .endofpacket
		.pixel_fondo               (avalon_st_adapter_001_out_0_data),                          //         background_sink.data
		.pixel_fondo_empty         (avalon_st_adapter_001_out_0_empty),                         //                        .empty
		.pixel_fondo_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),                   //                        .endofpacket
		.pixel_fondo_ready         (avalon_st_adapter_001_out_0_ready),                         //                        .ready
		.pixel_fondo_startofpacket (avalon_st_adapter_001_out_0_startofpacket),                 //                        .startofpacket
		.pixel_fondo_valid         (avalon_st_adapter_001_out_0_valid),                         //                        .valid
		.pixel_video               (avalon_st_adapter_002_out_0_data),                          //         foreground_sink.data
		.pixel_video_empty         (avalon_st_adapter_002_out_0_empty),                         //                        .empty
		.pixel_video_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),                   //                        .endofpacket
		.pixel_video_ready         (avalon_st_adapter_002_out_0_ready),                         //                        .ready
		.pixel_video_startofpacket (avalon_st_adapter_002_out_0_startofpacket),                 //                        .startofpacket
		.pixel_video_valid         (avalon_st_adapter_002_out_0_valid),                         //                        .valid
		.chipselect                (mm_interconnect_0_chromaprocessor_avalon_slave_chipselect), //            avalon_slave.chipselect
		.address                   (mm_interconnect_0_chromaprocessor_avalon_slave_address),    //                        .address
		.write                     (mm_interconnect_0_chromaprocessor_avalon_slave_write),      //                        .write
		.writedata                 (mm_interconnect_0_chromaprocessor_avalon_slave_writedata),  //                        .writedata
		.read                      (mm_interconnect_0_chromaprocessor_avalon_slave_read),       //                        .read
		.readdata                  (mm_interconnect_0_chromaprocessor_avalon_slave_readdata)    //                        .readdata
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (3),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_master_bfm (
		.clk                    (clk_50_in_clk),                  //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.avm_address            (mm_master_bfm_m0_address),       //        m0.address
		.avm_readdata           (mm_master_bfm_m0_readdata),      //          .readdata
		.avm_writedata          (mm_master_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest        (mm_master_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write              (mm_master_bfm_m0_write),         //          .write
		.avm_read               (mm_master_bfm_m0_read),          //          .read
		.avm_burstcount         (),                               // (terminated)
		.avm_begintransfer      (),                               // (terminated)
		.avm_beginbursttransfer (),                               // (terminated)
		.avm_byteenable         (),                               // (terminated)
		.avm_readdatavalid      (1'b0),                           // (terminated)
		.avm_arbiterlock        (),                               // (terminated)
		.avm_lock               (),                               // (terminated)
		.avm_debugaccess        (),                               // (terminated)
		.avm_transactionid      (),                               // (terminated)
		.avm_readid             (8'b00000000),                    // (terminated)
		.avm_writeid            (8'b00000000),                    // (terminated)
		.avm_clken              (),                               // (terminated)
		.avm_response           (2'b00),                          // (terminated)
		.avm_writeresponsevalid (1'b0),                           // (terminated)
		.avm_readresponse       (8'b00000000),                    // (terminated)
		.avm_writeresponse      (8'b00000000)                     // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (10),
		.ST_NUMSYMBOLS    (3),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (1),
		.VHDL_ID          (0)
	) st_sink_bfm (
		.clk                (clk_50_in_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_data          (avalon_st_adapter_out_0_data),          //      sink.data
		.sink_valid         (avalon_st_adapter_out_0_valid),         //          .valid
		.sink_ready         (avalon_st_adapter_out_0_ready),         //          .ready
		.sink_startofpacket (avalon_st_adapter_out_0_startofpacket), //          .startofpacket
		.sink_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //          .endofpacket
		.sink_empty         (2'b00),                                 // (terminated)
		.sink_channel       (1'b0),                                  // (terminated)
		.sink_error         (1'b0)                                   // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (10),
		.ST_NUMSYMBOLS    (3),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (1),
		.VHDL_ID          (0)
	) st_source_bfm_background (
		.clk               (clk_50_in_clk),                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),             // clk_reset.reset
		.src_data          (st_source_bfm_background_src_data),          //       src.data
		.src_valid         (st_source_bfm_background_src_valid),         //          .valid
		.src_ready         (st_source_bfm_background_src_ready),         //          .ready
		.src_startofpacket (st_source_bfm_background_src_startofpacket), //          .startofpacket
		.src_endofpacket   (st_source_bfm_background_src_endofpacket),   //          .endofpacket
		.src_empty         (),                                           // (terminated)
		.src_channel       (),                                           // (terminated)
		.src_error         ()                                            // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (10),
		.ST_NUMSYMBOLS    (3),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (1),
		.VHDL_ID          (0)
	) st_source_bfm_foreground (
		.clk               (clk_50_in_clk),                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),             // clk_reset.reset
		.src_data          (st_source_bfm_foreground_src_data),          //       src.data
		.src_valid         (st_source_bfm_foreground_src_valid),         //          .valid
		.src_ready         (st_source_bfm_foreground_src_ready),         //          .ready
		.src_startofpacket (st_source_bfm_foreground_src_startofpacket), //          .startofpacket
		.src_endofpacket   (st_source_bfm_foreground_src_endofpacket),   //          .endofpacket
		.src_empty         (),                                           // (terminated)
		.src_channel       (),                                           // (terminated)
		.src_error         ()                                            // (terminated)
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                      (clk_50_in_clk),                                             //                                    clk_50_clk.clk
		.mm_master_bfm_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // mm_master_bfm_clk_reset_reset_bridge_in_reset.reset
		.mm_master_bfm_m0_address                            (mm_master_bfm_m0_address),                                  //                              mm_master_bfm_m0.address
		.mm_master_bfm_m0_waitrequest                        (mm_master_bfm_m0_waitrequest),                              //                                              .waitrequest
		.mm_master_bfm_m0_read                               (mm_master_bfm_m0_read),                                     //                                              .read
		.mm_master_bfm_m0_readdata                           (mm_master_bfm_m0_readdata),                                 //                                              .readdata
		.mm_master_bfm_m0_write                              (mm_master_bfm_m0_write),                                    //                                              .write
		.mm_master_bfm_m0_writedata                          (mm_master_bfm_m0_writedata),                                //                                              .writedata
		.ChromaProcessor_avalon_slave_address                (mm_interconnect_0_chromaprocessor_avalon_slave_address),    //                  ChromaProcessor_avalon_slave.address
		.ChromaProcessor_avalon_slave_write                  (mm_interconnect_0_chromaprocessor_avalon_slave_write),      //                                              .write
		.ChromaProcessor_avalon_slave_read                   (mm_interconnect_0_chromaprocessor_avalon_slave_read),       //                                              .read
		.ChromaProcessor_avalon_slave_readdata               (mm_interconnect_0_chromaprocessor_avalon_slave_readdata),   //                                              .readdata
		.ChromaProcessor_avalon_slave_writedata              (mm_interconnect_0_chromaprocessor_avalon_slave_writedata),  //                                              .writedata
		.ChromaProcessor_avalon_slave_chipselect             (mm_interconnect_0_chromaprocessor_avalon_slave_chipselect)  //                                              .chipselect
	);

	nios_system_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_50_in_clk),                                         // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                        // in_rst_0.reset
		.in_0_data           (chromaprocessor_avalon_streaming_source_data),          //     in_0.data
		.in_0_valid          (chromaprocessor_avalon_streaming_source_valid),         //         .valid
		.in_0_ready          (chromaprocessor_avalon_streaming_source_ready),         //         .ready
		.in_0_startofpacket  (chromaprocessor_avalon_streaming_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (chromaprocessor_avalon_streaming_source_endofpacket),   //         .endofpacket
		.in_0_empty          (chromaprocessor_avalon_streaming_source_empty),         //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),                          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                 //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                    //         .endofpacket
	);

	nios_system_avalon_st_adapter_001 #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_50_in_clk),                              // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),             // in_rst_0.reset
		.in_0_data           (st_source_bfm_background_src_data),          //     in_0.data
		.in_0_valid          (st_source_bfm_background_src_valid),         //         .valid
		.in_0_ready          (st_source_bfm_background_src_ready),         //         .ready
		.in_0_startofpacket  (st_source_bfm_background_src_startofpacket), //         .startofpacket
		.in_0_endofpacket    (st_source_bfm_background_src_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),           //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),          //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),          //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket),  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),    //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)           //         .empty
	);

	nios_system_avalon_st_adapter_001 #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_002 (
		.in_clk_0_clk        (clk_50_in_clk),                              // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),             // in_rst_0.reset
		.in_0_data           (st_source_bfm_foreground_src_data),          //     in_0.data
		.in_0_valid          (st_source_bfm_foreground_src_valid),         //         .valid
		.in_0_ready          (st_source_bfm_foreground_src_ready),         //         .ready
		.in_0_startofpacket  (st_source_bfm_foreground_src_startofpacket), //         .startofpacket
		.in_0_endofpacket    (st_source_bfm_foreground_src_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_002_out_0_data),           //    out_0.data
		.out_0_valid         (avalon_st_adapter_002_out_0_valid),          //         .valid
		.out_0_ready         (avalon_st_adapter_002_out_0_ready),          //         .ready
		.out_0_startofpacket (avalon_st_adapter_002_out_0_startofpacket),  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),    //         .endofpacket
		.out_0_empty         (avalon_st_adapter_002_out_0_empty)           //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_50_in_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
